LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
--USE IEEE.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;
use IEEE.numeric_std.ALL;

ENTITY tb_placa IS
	PORT (CLOCK_50 : IN std_logic;
			SD_CLK  : OUT std_logic; -- sclk 
			SD_CMD  : OUT std_logic; -- mosi
			SD_DAT  : IN  std_logic; -- miso
			SD_DAT3 : OUT std_logic; -- ss_n
			
			SW   : IN std_logic_vector(9  DOWNTO 0);
			KEY  : IN std_logic_vector(0  DOWNTO 0);
			LEDR : OUT std_logic_vector(4 DOWNTO 0);
			
			HEX0 : OUT std_logic_vector(6 DOWNTO 0);
			HEX1 : OUT std_logic_vector(6 DOWNTO 0);
			HEX2 : OUT std_logic_vector(6 DOWNTO 0);
			HEX3 : OUT std_logic_vector(6 DOWNTO 0)
	);
END tb_placa;

ARCHITECTURE Structure OF tb_placa IS 

COMPONENT sd_controller is
generic (
	clockRate : integer := 50000000;		-- Incoming clock is 50MHz (can change this to 2000 to test Write Timeout)
	slowClockDivider : integer := 64;	-- Basic clock is 25MHz, slow clock for startup is 25/64 = 390kHz
	R1_TIMEOUT : integer := 10;			-- Number of bytes to wait before giving up on receiving R1 response
	WRITE_TIMEOUT : integer range 0 to 999 := 500		-- Number of ms to wait before giving up on write completing
	);
port (
	cs : out std_logic;				-- To SD card
	mosi : out std_logic;			-- To SD card
	miso : in std_logic;			-- From SD card
	sclk : out std_logic;			-- To SD card
	card_present : in std_logic;	-- From socket - can be fixed to '1' if no switch is present
	card_write_prot : in std_logic;	-- From socket - can be fixed to '0' if no switch is present, or '1' to make a Read-Only interface

	rd : in std_logic;				-- Trigger single block read
	-- rd_multiple : in std_logic;		-- Trigger multiple block read
	dout : out std_logic_vector(7 downto 0);	-- Data from SD card
	dout_avail : out std_logic;		-- Set when dout is valid
	dout_taken : in std_logic;		-- Acknowledgement for dout
	
	-- wr : in std_logic;				-- Trigger single block write
	-- wr_multiple : in std_logic;		-- Trigger multiple block write
	-- din : in std_logic_vector(7 downto 0);	-- Data to SD card
	-- din_valid : in std_logic;		-- Set when din is valid
	-- din_taken : out std_logic;		-- Ackowledgement for din
	
	addr : in std_logic_vector(31 downto 0);	-- Block address
	-- erase_count : in std_logic_vector(7 downto 0); -- For wr_multiple only

	sd_error : out std_logic;		-- '1' if an error occurs, reset on next RD or WR
	sd_busy : out std_logic;		-- '0' if a RD or WR can be accepted
	sd_error_code : out std_logic_vector(2 downto 0); -- See above, 000=No error
	
	
	reset : in std_logic;	-- System reset
	clk : in std_logic		-- twice the SPI clk (max 50MHz)
);
END COMPONENT;

COMPONENT sd_driver IS
    PORT ( addr  : IN std_logic_vector(15 downto 0);
			  rd    : IN std_logic;
			  busy : IN std_logic;
			  dout  : IN std_logic_vector(7 downto 0);
			  dout_avail : IN std_logic;
			  dout_taken : OUT std_logic;
			  data  : OUT std_logic_vector(15 downto 0) := (others => '0');
			  valid : OUT std_logic
);
END COMPONENT;

COMPONENT driverHex IS
	PORT (
		num : IN std_logic_vector(15 DOWNTO 0);
		display_en : IN std_logic_vector(3 downto 0);
		HEX0 : OUT std_logic_vector(6 DOWNTO 0);
		HEX1 : OUT std_logic_vector(6 DOWNTO 0);
		HEX2 : OUT std_logic_vector(6 DOWNTO 0);
		HEX3 : OUT std_logic_vector(6 DOWNTO 0)
	);
END COMPONENT;

signal reset : std_logic;

signal rd       : std_logic;
signal rd_debug : std_logic;
signal addr  : std_logic_vector(31 downto 0);
signal data  : std_logic_vector(15 downto 0);
signal valid : std_logic;

signal sd_busy    : std_logic;
signal dout       : std_logic_vector(7 downto 0);
signal dout_avail : std_logic;
signal dout_taken : std_logic;
signal cs         : std_logic;

signal sd_error      : std_logic;
signal sd_error_code : std_logic_vector(2 downto 0);

BEGIN

	SD_DAT3 <= not cs;
	rd <= '0' when SW(9) = '1'  else
			'1' when KEY(0) = '0' else 
					'0' when valid = '1'  else
					rd;
	LEDR(2) <= rd;
	LEDR(3) <= valid;
	--rd  <= rd_debug;
	reset   <= SW(9);
	addr    <= x"0000" & "0000000" & SW(8 downto 0);
	
	LEDR(0) <= valid;
	LEDR(1) <= sd_busy;
	
asdf: driverHex PORT MAP (
		num => data,
		display_en => "1111",
		HEX0 => HEX0,
		HEX1 => HEX1,
		HEX2 => HEX2,
		HEX3 => HEX3
	);

	-- Instantiate the Unit Under Test (UUT)
   uut: sd_controller PORT MAP (
          cs => cs,
          mosi => SD_CMD,
          miso => SD_DAT,
          sclk => SD_CLK,
			 card_present => '1',
			 card_write_prot => '0',
          -- sd_type => sd_state,
          -- sd_fsm => sd_fsm,
			 sd_error => sd_error,
			 sd_error_code => sd_error_code,
			 sd_busy => sd_busy,
          rd => rd,
          -- rd_multiple => rd_multiple,
          -- wr => wr,
          -- wr_multiple => wr_multiple,
          addr => addr,
			 -- erase_count => "00000010",
          reset => reset,
          -- din => din,
          -- din_valid => din_valid,
          -- din_taken => din_taken,
          dout => dout,
          dout_avail => dout_avail,
          dout_taken => dout_taken,
          clk => CLOCK_50
        );
		sd_drv: sd_driver PORT MAP (addr  => addr(15 downto 0),
																rd => rd,
																busy => sd_busy,
																dout => dout,
																dout_avail => dout_avail,
																dout_taken => dout_taken,
																data  => data,
																valid => valid);

END Structure;